module serial_paralelo1( output reg [7:0] data_rx000,
			 output reg valid_rx000, active,
			 input wire data_out, reset,
			 input wire clk_4f, clk_32f );

   // ESTRUCTURA DE ENTRADAS Y SALIDAS QUE SE DEBEN USAR
   // PARA QUE EXISTA COERENCIA
   
endmodule // serial_paralelo1

   
 

   
