module serial_paralelo2( output reg IDLE_OUT,
			 input wire clk_f, clk_4f, clk_32f,
			 input wire reset, inserter );

 // AL FINAL IDLE_OUT DEBE ESTAR SINCRONIZADO AL FLANCO ALTO clk_f

   
   
endmodule // serial_paralelo2

      
      
      
   
